CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 70 1680 1020
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 70 1680 1020
144179218 0
0
6 Title:
5 Name:
0
0
0
38
7 Ground~
168 243 209 0 1 3
0 0
0
0 0 53344 0
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 66 431 0 1 3
0 0
0
0 0 53344 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 240 597 0 1 3
0 0
0
0 0 53344 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
9 V Source~
197 239 565 0 1 5
0 0
0
0 0 17248 0
3 10V
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
6153 0 0
0
0
11 Signal Gen~
195 34 380 0 19 64
0 0 0 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
5 -1/1V
-18 -30 17 -22
2 V3
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
11 Signal Gen~
195 195 179 0 19 64
0 0 0 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
5 -1/1V
-18 -30 17 -22
2 V2
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
7734 0 0
0
0
9 Resistor~
219 280 529 0 1 5
0 0
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
7 Ground~
168 113 785 0 1 3
0 0
0
0 0 53344 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3747 0 0
0
0
2 +V
167 149 785 0 1 3
0 0
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3549 0 0
0
0
6 AD624~
219 252 748 0 1 25
0 0
0
0 0 4928 0
5 AD624
-18 -45 17 -37
2 U1
-7 -55 7 -47
0
0
44 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %10 %11 %12 %S
0
0
5 DIP16
25

0 16 1 2 7 6 9 8 3 10
13 12 11 16 1 2 7 6 9 8
3 10 13 12 11 0
88 0 0 256 1 0 0 0
1 U
7931 0 0
0
0
7 Ground~
168 264 437 0 1 3
0 0
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9325 0 0
0
0
9 Resistor~
219 229 421 0 1 5
0 0
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
10 Capacitor~
219 151 433 0 1 5
0 0
0
0 0 832 0
3 1uF
-11 -18 10 -10
3 C12
-11 -28 10 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3834 0 0
0
0
9 Resistor~
219 149 411 0 1 5
0 0
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 149 311 0 1 5
0 0
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
7 Ground~
168 503 537 0 1 3
0 0
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4718 0 0
0
0
7 Ground~
168 419 589 0 1 3
0 0
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3874 0 0
0
0
7 Ground~
168 324 586 0 1 3
0 0
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6671 0 0
0
0
7 Ground~
168 404 422 0 1 3
0 0
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3789 0 0
0
0
7 Ground~
168 325 420 0 1 3
0 0
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4871 0 0
0
0
7 Ground~
168 386 226 0 1 3
0 0
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3750 0 0
0
0
7 Ground~
168 318 225 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8778 0 0
0
0
10 Capacitor~
219 324 558 0 1 5
0 0
0
0 0 832 90
3 1uF
11 0 32 8
3 C11
11 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
538 0 0
0
0
10 Capacitor~
219 419 558 0 1 5
0 0
0
0 0 832 90
3 1uF
11 0 32 8
3 C10
11 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6843 0 0
0
0
9 Inductor~
219 369 529 0 1 5
0 0
0
0 0 832 0
3 1uH
-11 -17 10 -9
2 L4
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3136 0 0
0
0
10 Capacitor~
219 324 392 0 1 5
0 0
0
0 0 832 90
3 1uF
11 0 32 8
2 C9
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5950 0 0
0
0
10 Capacitor~
219 403 392 0 1 5
0 0
0
0 0 832 90
3 1uF
11 0 32 8
2 C8
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5670 0 0
0
0
10 Capacitor~
219 432 359 0 1 5
0 0
0
0 0 832 0
3 1uF
-11 -18 10 -10
2 C7
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6828 0 0
0
0
10 Capacitor~
219 291 357 0 1 5
0 0
0
0 0 832 0
3 1uF
-11 -18 10 -10
2 C6
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6735 0 0
0
0
9 Inductor~
219 364 358 0 1 5
0 0
0
0 0 832 0
3 1uH
-11 -17 10 -9
2 L3
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
8365 0 0
0
0
10 Capacitor~
219 288 174 0 1 5
0 0
0
0 0 832 0
3 1uF
-11 -18 10 -10
2 C5
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4132 0 0
0
0
10 Capacitor~
219 431 175 0 1 5
0 0
0
0 0 832 0
3 1uF
-11 -18 10 -10
2 C4
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4551 0 0
0
0
10 Capacitor~
219 319 196 0 1 5
0 0
0
0 0 832 90
3 1uF
11 0 32 8
2 C3
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3635 0 0
0
0
10 Capacitor~
219 386 197 0 1 5
0 0
0
0 0 832 90
3 1uF
11 0 32 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3973 0 0
0
0
9 Inductor~
219 355 176 0 1 5
0 0
0
0 0 832 0
3 1uH
-11 -17 10 -9
2 L2
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3851 0 0
0
0
10 Capacitor~
219 818 334 0 1 5
0 0
0
0 0 832 90
3 1uF
11 0 32 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8383 0 0
0
0
9 Resistor~
219 861 352 0 1 5
0 0
0
0 0 864 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9334 0 0
0
0
9 Inductor~
219 861 317 0 1 5
0 0
0
0 0 832 270
3 1uH
6 -4 27 4
2 L1
10 -14 24 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
7471 0 0
0
0
43
1 1 0 0 0 0 0 6 31 0 0 2
226 174
279 174
2 1 0 0 0 0 0 6 1 0 0 3
226 184
243 184
243 203
1 0 0 0 0 0 0 5 0 0 17 2
65 375
80 375
2 1 0 0 0 0 0 5 2 0 0 3
65 385
66 385
66 425
2 1 0 0 0 0 0 4 3 0 0 3
239 586
240 586
240 591
1 1 0 0 0 0 0 4 7 0 0 3
239 544
239 529
262 529
0 5 0 0 0 0 0 0 10 8 0 5
309 529
309 676
183 676
183 748
219 748
2 0 0 0 0 0 0 7 0 0 26 2
298 529
324 529
1 7 0 0 0 0 0 9 10 0 0 3
149 794
219 794
219 766
8 10 0 0 0 0 0 10 10 0 0 6
219 739
211 739
211 685
296 685
296 730
285 730
4 1 0 0 0 0 0 10 8 0 0 3
219 757
113 757
113 779
3 0 0 0 0 0 0 10 0 0 16 3
219 721
199 721
199 311
0 2 0 0 0 0 0 0 10 18 0 3
192 421
192 730
219 730
9 6 0 0 0 0 0 10 10 0 0 2
285 757
285 766
2 1 0 0 0 0 0 12 11 0 0 3
247 421
264 421
264 431
2 1 0 0 0 0 0 15 29 0 0 4
167 311
267 311
267 357
282 357
1 0 0 0 0 0 0 15 0 0 20 4
131 311
80 311
80 423
113 423
1 0 0 0 0 0 0 12 0 0 19 2
211 421
176 421
2 2 0 0 0 0 0 13 14 0 0 4
160 433
176 433
176 411
167 411
1 1 0 0 0 0 0 14 13 0 0 4
131 411
113 411
113 433
142 433
0 0 0 0 0 0 0 0 0 23 42 3
469 266
845 266
845 293
2 0 0 0 0 0 0 28 0 0 23 2
441 359
469 359
0 2 0 0 0 0 0 0 32 25 0 4
419 529
469 529
469 175
440 175
0 1 0 0 0 0 0 0 16 41 0 4
845 382
845 501
503 501
503 531
2 2 0 0 0 0 0 25 24 0 0 3
387 529
419 529
419 549
2 1 0 0 0 0 0 23 25 0 0 3
324 549
324 529
351 529
1 1 0 0 0 0 0 17 24 0 0 2
419 583
419 567
1 1 0 0 0 0 0 18 23 0 0 2
324 580
324 567
1 1 0 0 0 0 0 27 19 0 0 3
403 401
404 401
404 416
1 1 0 0 0 0 0 26 20 0 0 3
324 401
325 401
325 414
2 0 0 0 0 0 0 26 0 0 34 2
324 383
324 358
2 0 0 0 0 0 0 27 0 0 33 2
403 383
403 359
2 1 0 0 0 0 0 30 28 0 0 3
382 358
382 359
423 359
2 1 0 0 0 0 0 29 30 0 0 3
300 357
300 358
346 358
1 1 0 0 0 0 0 33 22 0 0 3
319 205
318 205
318 219
1 1 0 0 0 0 0 34 21 0 0 2
386 206
386 220
2 0 0 0 0 0 0 34 0 0 39 2
386 188
386 175
0 2 0 0 0 0 0 0 33 40 0 2
319 176
319 187
2 1 0 0 0 0 0 35 32 0 0 3
373 176
373 175
422 175
2 1 0 0 0 0 0 31 35 0 0 3
297 174
297 176
337 176
1 1 0 0 0 0 0 37 36 0 0 4
861 370
861 382
818 382
818 343
2 1 0 0 0 0 0 36 38 0 0 4
818 325
818 293
861 293
861 299
2 2 0 0 0 0 0 37 38 0 0 2
861 334
861 335
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
